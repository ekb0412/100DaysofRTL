`timescale 1ns / 1ps

module tb_nor;
    reg a, b;
    wire nor_out;
         
    decoder_nor dut(a, b, nor_out);
    initial begin
            a= 1'b0; b= 1'b0;
        #10 a= 1'b0; b= 1'b1;
        #10 a= 1'b1; b= 1'b0;
        #10 a= 1'b1; b= 1'b1;
    end
    initial 
     begin $monitor("a: %b  b: %b  nor: %b ",a, b, nor_out);
     #40 $finish;
     end
endmodule
